

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO spc2 
  PIN Cfg_in 
    ANTENNAPARTIALMETALAREA 2.6656 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.1392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.198 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.9359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 133.646 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.791919 LAYER V3 ;
  END Cfg_in
  PIN Clk 
    ANTENNAPARTIALMETALAREA 26.3424 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2534 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.7539 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 150.975 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.58384 LAYER V3 ;
  END Clk
  PIN Resetn 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 6.3504 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.0416 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 14.652 LAYER M4 ; 
    ANTENNAMAXAREACAR 16.2465 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 57.0702 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.79727 LAYER V4 ;
  END Resetn
  PIN F[3] 
    ANTENNADIFFAREA 0.9488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.784 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.688 LAYER M3 ;
  END F[3]
  PIN F[2] 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.0368 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.9664 LAYER M4 ;
  END F[2]
  PIN F[1] 
    ANTENNADIFFAREA 0.9488 LAYER M3 ; 
  END F[1]
  PIN F[0] 
    ANTENNADIFFAREA 0.9488 LAYER M3 ; 
  END F[0]
  PIN IQ 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.1136 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 34.944 LAYER M4 ;
  END IQ
  PIN GS[3] 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 12.152 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.9328 LAYER M4 ;
  END GS[3]
  PIN GS[2] 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.2912 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.2672 LAYER M4 ;
  END GS[2]
  PIN GS[1] 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.4688 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.5904 LAYER M4 ;
  END GS[1]
  PIN GS[0] 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.312 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.0528 LAYER M4 ;
  END GS[0]
  PIN CE 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.7232 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8912 LAYER M4 ;
  END CE
  PIN NS 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.4688 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.5904 LAYER M4 ;
  END NS
  PIN GD[2] 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.4288 LAYER M4 ;
  END GD[2]
  PIN GD[1] 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.1136 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 34.944 LAYER M4 ;
  END GD[1]
  PIN GD[0] 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.7024 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.1056 LAYER M4 ;
  END GD[0]
  PIN FS 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.9488 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.4688 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.5904 LAYER M4 ;
  END FS
  PIN RE 
    ANTENNADIFFAREA 0.9488 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.624 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.568 LAYER M3 ;
  END RE
END spc2

END LIBRARY
