/*
 * Hello World for Papillio Duo
 * Author: Saul Rodriguez
 * Date: 2016-09-09
 *
 */
 
 module hello(in,out);
 
 input in;
 output out;
 
 assign out = ~in;
  
 endmodule 
 
 
