

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO sar5 
  PIN clk 
    ANTENNAPARTIALMETALAREA 26.6168 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.7952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.584 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.2015 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 105.688 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38586 LAYER V3 ;
  END clk
  PIN comp 
    ANTENNAPARTIALMETALAREA 15.9992 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 54.8544 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8032 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.423 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.0912 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.327 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.9596 LAYER V3 ;
  END comp
  PIN resetn 
    ANTENNAPARTIALMETALAREA 17.0968 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 58.6176 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.168 LAYER M4 ; 
    ANTENNAMAXAREACAR 13.0543 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 45.1121 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.346465 LAYER V4 ;
  END resetn
  PIN out[4] 
    ANTENNADIFFAREA 1.442 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 15.9544 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.7008 LAYER M3 ;
  END out[4]
  PIN out[3] 
    ANTENNADIFFAREA 1.127 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.1176 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 48.4032 LAYER M2 ;
  END out[3]
  PIN out[2] 
    ANTENNADIFFAREA 1.442 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.4 LAYER M2 ;
  END out[2]
  PIN out[1] 
    ANTENNADIFFAREA 1.442 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 14.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.4 LAYER M2 ;
  END out[1]
  PIN out[0] 
    ANTENNADIFFAREA 1.442 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.3864 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.3248 LAYER M3 ;
  END out[0]
END sar5

END LIBRARY
