

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO nnspc 
  PIN Cfg_in 
    ANTENNAPARTIALMETALAREA 2.352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.198 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.6106 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 178.73 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.58384 LAYER V3 ;
  END Cfg_in
  PIN Clk 
    ANTENNAPARTIALMETALAREA 2.8616 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.08 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.269 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.99648 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 21.2753 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.858238 LAYER V3 ;
  END Clk
  PIN Resetn 
    ANTENNAPARTIALMETALAREA 0.1568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5376 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2196 LAYER M3 ; 
    ANTENNAMAXAREACAR 23.0647 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 81.1776 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.42805 LAYER V3 ;
  END Resetn
  PIN NSEL[4] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 1.274 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.0544 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.1696 LAYER M4 ;
  END NSEL[4]
  PIN NSEL[3] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 1.274 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.5248 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.7824 LAYER M4 ;
  END NSEL[3]
  PIN NSEL[2] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 1.274 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.4272 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.0192 LAYER M4 ;
  END NSEL[2]
  PIN NSEL[1] 
    ANTENNADIFFAREA 1.274 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.9128 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.1296 LAYER M3 ;
  END NSEL[1]
  PIN NSEL[0] 
    ANTENNAPARTIALMETALAREA 0.308 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 1.274 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.1936 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.504 LAYER M4 ;
  END NSEL[0]
  PIN DAC[3] 
    ANTENNAPARTIALMETALAREA 0.188 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 1.274 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.232 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.4928 LAYER M4 ;
  END DAC[3]
  PIN DAC[2] 
    ANTENNADIFFAREA 1.274 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.9336 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9152 LAYER M3 ;
  END DAC[2]
  PIN DAC[1] 
    ANTENNADIFFAREA 1.274 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.3272 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5504 LAYER M3 ;
  END DAC[1]
  PIN DAC[0] 
    ANTENNADIFFAREA 1.274 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.2088 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0016 LAYER M3 ;
  END DAC[0]
  PIN RE 
    ANTENNADIFFAREA 1.274 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.6184 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.0048 LAYER M3 ;
  END RE
END nnspc

END LIBRARY
