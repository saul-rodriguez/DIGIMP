/**************************************
* Module: spc2
* Date:2015-11-08  
* Author: saul     
*
* Description: Serial to Parallel converter used for configuring BIO IC V1
* This block uses 3 control lines: Cfg_in, Clk, and Resetn 
* Cfg_in is sampled at rising edge of Clk. After 14 bits, the data is latched to the paralell outputs
* 
* 
* Configuation word: F3,F2,F1,F0,    IQ,   GS3,GS2,GS1,GS0,  CE,   NS,    GD2,GD1,GD0
* F<3:0>    Frequency selection 0 - 15  (0 highest frequency (VCO freq), 15 lowest frequency)
* IQ        I = 0, Q = 1
* GS<3:0>   Signal Generator Gain [0000, 0001, 0011, 0111, 1111]
* CE        Signal Generator enable 
* NS        Signal Generator number of steps NS = 0 (32 steps), NS = 1 (16 steps)
* GD<2:0>   Demodulator Gain [100, 101, 111, 011] (NOTE: G[2] is active low logic!)
* FS        Filter Selection FS = 0 (fast), FS = 1 (slow)
* RE        Reserve pin
* 
***************************************/
module  spc2(
Cfg_in,
Clk,
Resetn,
F,
IQ,
GS,
CE,
NS,
GD,
FS,
RE
);

input Cfg_in, Clk, Resetn;

output reg[3:0] F;
output reg IQ;
output reg [3:0] GS;
output reg CE;
output reg NS;
output reg [2:0] GD;
output reg FS;
output reg RE;

reg [15:0] out; 
reg [4:0] count;

wire strobe;

/*
* Right Shift register with async. reset  
*/
always @(posedge Clk, negedge Resetn)
begin
    if (Resetn == 0) begin
        out <= 0;
        count <= 16;
    end else begin
        //Shift the data
        out[15] <= Cfg_in;
        out[14] <= out[15];
        out[13] <= out[14];
        out[12] <= out[13];
        out[11] <= out[12];
        out[10] <= out[11];
        out[9] <= out[10];
        out[8] <= out[9];
        out[7] <= out[8];
        out[6] <= out[7];
        out[5] <= out[6];
        out[4] <= out[5];
        out[3] <= out[4];
        out[2] <= out[3];
        out[1] <= out[2];
        out[0] <= out[1];
        
        //Decrement the counter
        count <= count - 1;
    end    
end

assign strobe = (!count) & (~Clk);

always @(posedge strobe, negedge Resetn)
begin
    if (Resetn == 0) begin
        F[3:0] <= 0;
        IQ <= 0;
        GS[3:0] <= 0;
        CE <= 0;
        NS <= 0;
        GD[2:0] <= 0;
        FS <= 0;
        RE <= 0;
    end else begin
        F[3:0] <= out[15:12];
        IQ <= out[11];
        GS[3:0] <= out[10:7];
        CE <= out[6];
        NS <= out[5];
        GD[2:0] <= out[4:2];
        FS <= out[1];
        RE <= out[0];
    end
end

endmodule











