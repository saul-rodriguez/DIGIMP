

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO fet_dec 
  PIN in[4] 
    ANTENNAPARTIALMETALAREA 3.9984 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.9776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6912 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.7481 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.901 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.9596 LAYER V3 ;
  END in[4]
  PIN in[3] 
    ANTENNAPARTIALMETALAREA 0.1176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 8.0752 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9552 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3852 LAYER M4 ; 
    ANTENNAMAXAREACAR 45.0477 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 160.061 LAYER M4 ;
    ANTENNAMAXCUTCAR 2.79392 LAYER V4 ;
  END in[3]
  PIN in[2] 
    ANTENNAPARTIALMETALAREA 1.6856 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.7792 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4068 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.998 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 94.9031 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.36525 LAYER V3 ;
  END in[2]
  PIN in[1] 
    ANTENNAPARTIALMETALAREA 9.4472 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.1968 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6552 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.0708 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 218.352 LAYER M3 ;
    ANTENNAMAXCUTCAR 4.93082 LAYER V3 ;
  END in[1]
  PIN in[0] 
    ANTENNAPARTIALMETALAREA 8.7024 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.1056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5256 LAYER M3 ; 
    ANTENNAMAXAREACAR 57.2695 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 199.851 LAYER M3 ;
    ANTENNAMAXCUTCAR 3.07451 LAYER V3 ;
  END in[0]
  PIN out[31] 
    ANTENNAPARTIALMETALAREA 0.2352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.7056 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.688 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V4 ;
    ANTENNADIFFAREA 1.2688 LAYER MT ; 
    ANTENNAPARTIALMETALAREA 11.6816 LAYER MT ;
    ANTENNAPARTIALMETALSIDEAREA 40.32 LAYER MT ;
  END out[31]
  PIN out[30] 
    ANTENNAPARTIALMETALAREA 0.1176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.9952 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.3952 LAYER M4 ;
  END out[30]
  PIN out[29] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.1168 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5264 LAYER M3 ;
  END out[29]
  PIN out[28] 
    ANTENNAPARTIALMETALAREA 0.2352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.1328 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 38.7072 LAYER M4 ;
  END out[28]
  PIN out[27] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.1568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5376 LAYER M3 ;
  END out[27]
  PIN out[26] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.0576 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.752 LAYER M3 ;
  END out[26]
  PIN out[25] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.1152 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.504 LAYER M3 ;
  END out[25]
  PIN out[24] 
    ANTENNAPARTIALMETALAREA 0.1568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5376 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.2704 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 35.4816 LAYER M4 ;
  END out[24]
  PIN out[23] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.2136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.144 LAYER M3 ;
  END out[23]
  PIN out[22] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.9888 LAYER M3 ;
  END out[22]
  PIN out[21] 
    ANTENNAPARTIALMETALAREA 0.196 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.672 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 1.2688 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 13.2496 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.696 LAYER M4 ;
  END out[21]
  PIN out[20] 
    ANTENNAPARTIALMETALAREA 4.4688 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.5904 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.4304 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6016 LAYER M4 ;
  END out[20]
  PIN out[19] 
    ANTENNAPARTIALMETALAREA 0.1176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 1.2688 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 11.6032 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 40.32 LAYER M4 ;
  END out[19]
  PIN out[18] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.0752 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9552 LAYER M3 ;
  END out[18]
  PIN out[17] 
    ANTENNAPARTIALMETALAREA 0.2352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.3888 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 29.0304 LAYER M4 ;
  END out[17]
  PIN out[16] 
    ANTENNAPARTIALMETALAREA 0.2352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.7232 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8912 LAYER M4 ;
  END out[16]
  PIN out[15] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.7232 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8912 LAYER M3 ;
  END out[15]
  PIN out[14] 
    ANTENNAPARTIALMETALAREA 0.1568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5376 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.7408 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 37.0944 LAYER M4 ;
  END out[14]
  PIN out[13] 
    ANTENNAPARTIALMETALAREA 0.1568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5376 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 10.5056 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.5568 LAYER M4 ;
  END out[13]
  PIN out[12] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.1368 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1664 LAYER M3 ;
  END out[12]
  PIN out[11] 
    ANTENNAPARTIALMETALAREA 0.2352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9.016 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 31.1808 LAYER M4 ;
  END out[11]
  PIN out[10] 
    ANTENNAPARTIALMETALAREA 0.1176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 0.8624 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2256 LAYER M4 ;
  END out[10]
  PIN out[9] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.3712 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8272 LAYER M3 ;
  END out[9]
  PIN out[8] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.8976 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.632 LAYER M3 ;
  END out[8]
  PIN out[7] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.2912 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.2672 LAYER M3 ;
  END out[7]
  PIN out[6] 
    ANTENNAPARTIALMETALAREA 1.0192 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7632 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 7.2912 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.2672 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V4 ;
    ANTENNADIFFAREA 1.2688 LAYER MT ; 
    ANTENNAPARTIALMETALAREA 8.3888 LAYER MT ;
    ANTENNAPARTIALMETALSIDEAREA 29.0304 LAYER MT ;
  END out[6]
  PIN out[5] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.9008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.2144 LAYER M3 ;
  END out[5]
  PIN out[4] 
    ANTENNAPARTIALMETALAREA 0.1176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.0368 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.9664 LAYER M4 ;
  END out[4]
  PIN out[3] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.528 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3648 LAYER M3 ;
  END out[3]
  PIN out[2] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.2704 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.4816 LAYER M3 ;
  END out[2]
  PIN out[1] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.4896 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.376 LAYER M3 ;
  END out[1]
  PIN out[0] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.6272 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1504 LAYER M3 ;
  END out[0]
END fet_dec

END LIBRARY
