/**************************************
* Module: DacCtrl
* Date:2015-09-25  
* Author: saul     
*
* Description: 
* 
*  output P     32 steps    16 steps    8 step
* ------------------------------------------
* 8             1         1          1
* 7             0.9808      
* 6             0.9239    0.9239  
* 5             0.8315      
* 4             0.7071    0.7071     0.7071
* 3             0.5556      
* 2             0.3827    0.3827  
* 1             0.1951      
* 0             0         0          0
* 9             -0.1951     
* 10            -0.3827   -0.3827 
* 11            -0.5556     
* 12            -0.7071   -0.7071    -0.7071
* 13            -0.8315     
* 14            -0.9239   -0.9239 
* 15            -0.9808     
* 16            -1        -1         -1
* 
* The I/Q signals are ahead of the sinusoidal signal:
* 32 steps:1/32*1/2*360 = 5.625 deg
* 16 steps: = 1/16*1/2*360 = 11.25 deg
* 
***************************************/

module  DacCtrl(
CountEnable,
Clk,
Resetn,
StepNum,
P,
IP,
IN,
QP,
QN
);


//Inputs
input CountEnable;
input Clk;
input Resetn;
input StepNum;


//Outputs
//output wire P1,P2,P3,P4,P5; //Control signals for the DAC
output reg [16:0] P; //Control signals for the DAC
output reg IP; // in-phase (I) reference clock
output reg QP; // quadrature (Q) reference clock
//output wire QP; // quadrature (Q) reference clock
output wire IN,QN; 

reg [16:0] S32;
reg [16:0] S16;

reg [4:0] count;

reg aux_Q;

// 5bit counter state machine
always @(posedge Clk, negedge Resetn)
begin
    if (Resetn == 0) begin
        count <= 0;
    end else begin
        count <= count + 1;    
    end    
end

// AMS VERSION 32 steps - 16 steps

//Intermediate signals 32 steps
always @(CountEnable, count)
begin
    if (CountEnable == 1) begin
        case(count)
            0:  S32 = 17'b0_0000_0000_0000_0001; //0 0V                
            1:  S32 = 17'b0_0000_0000_0000_0010;
            2:  S32 = 17'b0_0000_0000_0000_0100;
            3:  S32 = 17'b0_0000_0000_0000_1000;
            4:  S32 = 17'b0_0000_0000_0001_0000;
            5:  S32 = 17'b0_0000_0000_0010_0000;
            6:  S32 = 17'b0_0000_0000_0100_0000;
            7:  S32 = 17'b0_0000_0000_1000_0000;
            8:  S32 = 17'b0_0000_0001_0000_0000; //8 +1V
            9:  S32 = 17'b0_0000_0000_1000_0000;
            10: S32 = 17'b0_0000_0000_0100_0000;
            11: S32 = 17'b0_0000_0000_0010_0000;
            12: S32 = 17'b0_0000_0000_0001_0000;
            13: S32 = 17'b0_0000_0000_0000_1000;
            14: S32 = 17'b0_0000_0000_0000_0100;
            15: S32 = 17'b0_0000_0000_0000_0010;
            16: S32 = 17'b0_0000_0000_0000_0001;// 0V
            17: S32 = 17'b0_0000_0010_0000_0000; 
            18: S32 = 17'b0_0000_0100_0000_0000;
            19: S32 = 17'b0_0000_1000_0000_0000;
            20: S32 = 17'b0_0001_0000_0000_0000;
            21: S32 = 17'b0_0010_0000_0000_0000;
            22: S32 = 17'b0_0100_0000_0000_0000;
            23: S32 = 17'b0_1000_0000_0000_0000;            
            24: S32 = 17'b1_0000_0000_0000_0000; //16 -1V
            25: S32 = 17'b0_1000_0000_0000_0000;
            26: S32 = 17'b0_0100_0000_0000_0000;
            27: S32 = 17'b0_0010_0000_0000_0000;
            28: S32 = 17'b0_0001_0000_0000_0000;
            29: S32 = 17'b0_0000_1000_0000_0000;
            30: S32 = 17'b0_0000_0100_0000_0000;
            31: S32 = 17'b0_0000_0010_0000_0000;
            default: S32 = 17'b0_0000_0000_0000_0001; //0 0V
         endcase   
         
    end else begin
            S32 = 17'b0_0000_0000_0000_0001; //0 0V  
    end
end

//Intermediate signals 16 steps
always @(CountEnable, count)
begin
    if (CountEnable == 1) begin
        case(count)
            0:  S16 = 17'b0_0000_0000_0000_0001; //0 0V                
            1:  S16 = 17'b0_0000_0000_0000_0100;
            2:  S16 = 17'b0_0000_0000_0001_0000;
            3:  S16 = 17'b0_0000_0000_0100_0000;
            4:  S16 = 17'b0_0000_0001_0000_0000;//8 +1V
            5:  S16 = 17'b0_0000_0000_0100_0000;
            6:  S16 = 17'b0_0000_0000_0001_0000;
            7:  S16 = 17'b0_0000_0000_0000_0100;
            8:  S16 = 17'b0_0000_0000_0000_0001; //0 0V
            9:  S16 = 17'b0_0000_0100_0000_0000;
            10: S16 = 17'b0_0001_0000_0000_0000;
            11: S16 = 17'b0_0100_0000_0000_0000;
            12: S16 = 17'b1_0000_0000_0000_0000; //16 -1V
            13: S16 = 17'b0_0100_0000_0000_0000;
            14: S16 = 17'b0_0001_0000_0000_0000;
            15: S16 = 17'b0_0000_0100_0000_0000;            
            16:  S16 = 17'b0_0000_0000_0000_0001; //0 0V                
            17:  S16 = 17'b0_0000_0000_0000_0100;
            18:  S16 = 17'b0_0000_0000_0001_0000;
            19:  S16 = 17'b0_0000_0000_0100_0000;
            20:  S16 = 17'b0_0000_0001_0000_0000;//8 +1V
            21:  S16 = 17'b0_0000_0000_0100_0000;
            22:  S16 = 17'b0_0000_0000_0001_0000;
            23:  S16 = 17'b0_0000_0000_0000_0100;
            24:  S16 = 17'b0_0000_0000_0000_0001; //0 0V
            25:  S16 = 17'b0_0000_0100_0000_0000;
            26: S16 = 17'b0_0001_0000_0000_0000;
            27: S16 = 17'b0_0100_0000_0000_0000;
            28: S16 = 17'b1_0000_0000_0000_0000; //16 -1V
            29: S16 = 17'b0_0100_0000_0000_0000;
            30: S16 = 17'b0_0001_0000_0000_0000;
            31: S16 = 17'b0_0000_0100_0000_0000;
                 
           
            default: S16 = 17'b0_0000_0000_0000_0001; //0 0V
         endcase   
         
    end else begin
            S16 = 17'b0_0000_0000_0000_0001; //0 0V  
    end
end

always @(StepNum,S16,S32)
begin
    if (StepNum == 0) begin // 0 selects 32 steps, 1 selects 16 steps
        P = S32;
    end else begin
        P = S16;
    end
    
end

// I/Q Outputs

always @(StepNum,count)
begin
    if(StepNum == 0) begin // 32 Steps
        IP <= ~count[4];
       
    end else begin // 16 steps
        IP <= ~count[3];
      
    end
end

assign IN = ~IP;


//Q is created by sampling I exactly in the middle of the high pulse. 
//Aux_Q is the clock used to sample I;
always @(StepNum,count)
begin
    if(StepNum == 0) begin //32 steps
        aux_Q = count[3];
    end else begin //16 steps
        aux_Q = count[2];
    end
end

always @(posedge aux_Q, negedge Resetn)
begin
    if (Resetn == 0) begin
        QP <= 0;         
    end else begin
        QP <= IP; 
    end    
end

assign QN = ~QP;

endmodule

