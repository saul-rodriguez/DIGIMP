

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO cur_dec 
  PIN out[15] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 10.1136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.944 LAYER M3 ;
  END out[15]
  PIN out[14] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 9.1728 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.7184 LAYER M3 ;
  END out[14]
  PIN out[13] 
    ANTENNAPARTIALMETALAREA 0.1176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.4096 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.816 LAYER M4 ;
  END out[13]
  PIN out[12] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 5.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.4288 LAYER M3 ;
  END out[12]
  PIN out[11] 
    ANTENNAPARTIALMETALAREA 0.1568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5376 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.88 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.4288 LAYER M4 ;
  END out[11]
  PIN out[10] 
    ANTENNAPARTIALMETALAREA 0.2352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.0752 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.9552 LAYER M4 ;
  END out[10]
  PIN out[9] 
    ANTENNAPARTIALMETALAREA 0.1176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.9184 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.4176 LAYER M4 ;
  END out[9]
  PIN out[8] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3008 LAYER M3 ;
  END out[8]
  PIN out[7] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.1568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5376 LAYER M3 ;
  END out[7]
  PIN out[6] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.6464 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9136 LAYER M3 ;
  END out[6]
  PIN out[5] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.8624 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2256 LAYER M3 ;
  END out[5]
  PIN out[4] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 3.528 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3648 LAYER M3 ;
  END out[4]
  PIN out[3] 
    ANTENNAPARTIALMETALAREA 0.1176 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4032 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.4304 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6016 LAYER M4 ;
  END out[3]
  PIN out[2] 
    ANTENNAPARTIALMETALAREA 0.2352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8064 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.9392 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2032 LAYER M4 ;
  END out[2]
  PIN out[1] 
    ANTENNAPARTIALMETALAREA 0.1568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5376 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNADIFFAREA 0.9464 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 7.6048 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 26.3424 LAYER M4 ;
  END out[1]
  PIN out[0] 
    ANTENNADIFFAREA 0.9464 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.252 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.1328 LAYER M3 ;
  END out[0]
  PIN in[3] 
    ANTENNAPARTIALMETALAREA 1.568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.376 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3852 LAYER M3 ; 
    ANTENNAMAXAREACAR 65.9183 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 239.519 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.38686 LAYER V3 ;
  END in[3]
  PIN in[2] 
    ANTENNAPARTIALMETALAREA 2.1168 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5264 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7848 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.0801 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 138.913 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.84886 LAYER V3 ;
  END in[2]
  PIN in[1] 
    ANTENNAPARTIALMETALAREA 3.9984 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.9776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4716 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.2678 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.829 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.65508 LAYER V3 ;
  END in[1]
  PIN in[0] 
    ANTENNAPARTIALMETALAREA 4.3904 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.0528 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.153 LAYER M3 ; 
    ANTENNAMAXAREACAR 58.1346 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 202.306 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER V3 ;
    ANTENNAMAXCUTCAR 3.07451 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 6.9776 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 24.192 LAYER M4 ;
    ANTENNAGATEAREA 0.5256 LAYER M4 ; 
    ANTENNAMAXAREACAR 71.4101 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 248.333 LAYER M4 ;
    ANTENNAMAXCUTCAR 3.07451 LAYER V4 ;
  END in[0]
END cur_dec

END LIBRARY
